module not_gate(y, a);
output y;
input a;

assign y = a;
endmodule
